module redict

interface Any {}
